library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
library work;
use work.dlxlib.all;

entity dlx_decode is
    Port ( 
        clk : in  STD_LOGIC;
        rst_l : in  STD_LOGIC := '0';
        addr_in : in STD_LOGIC_VECTOR (ADDR_WIDTH-1 downto 0);
        instr_in : in STD_LOGIC_VECTOR (INSTR_WIDTH-1 downto 0);
        writeback_data : in STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
        writeback_reg : in STD_LOGIC_VECTOR (4 downto 0);
        writeback_en : in STD_LOGIC;
        rs1_data : out STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
        rs2_data : out STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
        immediate : out STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);
        instr_out : out STD_LOGIC_VECTOR (INSTR_WIDTH-1 downto 0);
        addr_out : out STD_LOGIC_VECTOR (ADDR_WIDTH-1 downto 0)
    );
end dlx_decode;

architecture hierarchial of dlx_decode is

    signal opcode : STD_LOGIC_VECTOR (5 downto 0);
    signal rs1 : STD_LOGIC_VECTOR (4 downto 0);
    signal rs2 : STD_LOGIC_VECTOR (4 downto 0);
    signal imm16 : STD_LOGIC_VECTOR (15 downto 0);
    signal EX_instr : STD_LOGIC_VECTOR (INSTR_WIDTH-1 downto 0) := (others => '0');
    signal MEM_instr : STD_LOGIC_VECTOR (INSTR_WIDTH-1 downto 0) := (others => '0');
    signal WB_instr : STD_LOGIC_VECTOR (INSTR_WIDTH-1 downto 0) := (others => '0');

    component register_mem
        port (
            clk : in std_logic;
            read_addr1 : in std_logic_vector(4 downto 0);
            read_addr2 : in std_logic_vector(4 downto 0);
            write_addr : in std_logic_vector(4 downto 0);
            write_data : in std_logic_vector(DATA_WIDTH-1 downto 0);
            write_en : in std_logic := '0';
            read_q1 : out std_logic_vector(DATA_WIDTH-1 downto 0);
            read_q2 : out std_logic_vector(DATA_WIDTH-1 downto 0)
        );
    end component;

    component signExtend
        port ( 
            input : in  STD_LOGIC_VECTOR (15 downto 0);
            us : in STD_LOGIC;
            output : out  STD_LOGIC_VECTOR (31 downto 0)
        );
    end component;

    signal next_immediate : STD_LOGIC_VECTOR (DATA_WIDTH-1 downto 0);

begin

    opcode <= instr_in(31 downto 26);
    rs1 <= instr_in(20 downto 16);
    imm16 <= instr_in(15 downto 0);
    EX_instr <= instr_out;


    process(opcode) begin
        if opcode = SW then
            rs2 <= instr_in(25 downto 21);
        else
            rs2 <= instr_in(15 downto 11);
        end if;
    end process;

    register_inst : register_mem
        port map (
            clk => clk,
            read_addr1 => rs1,
            read_addr2 => rs2,
            write_addr => writeback_reg,
            write_data => writeback_data,
            write_en => writeback_en,
            read_q1 => rs1_data,
            read_q2 => rs2_data
        );

    signExtend_inst : signExtend
        port map (
            input => imm16,
            us => is_unsigned(opcode),
            output => next_immediate
        );


    process(clk, rst_l) begin
        if rising_edge(clk) then
            WB_instr <= MEM_instr;
            MEM_instr <= EX_instr;
            instr_out <= instr_in;
            addr_out <= addr_in;
            immediate <= next_immediate;
        end if;
    end process;

    process(instr_in, EX_instr, MEM_instr, WB_instr, rs1, rs2) begin
        if rs1 = EX_instr(25 downto 21) then
            
    end process;

end hierarchial;
