package dlxlib is
    constant ADDR_WIDTH : integer := 10;
    constant DATA_WIDTH : integer := 32;
    constant MEM_SIZE : integer := 2**ADDR_WIDTH;
end package dlxlib;