use IEEE.STD_LOGIC_1164.ALL;
use dlxlib.all;

entity mux is
    Parameter (
        N : integer := 2
        
    )