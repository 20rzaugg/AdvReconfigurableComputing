library IEEE;
use IEEE.std_logic_1164.all;

package LCM_PACKAGE is

    constant DATA_WIDTH : integer := 64;

end package LCM_PACKAGE;